CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
50
13 Logic Switch~
5 898 803 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21344 512
2 5V
-7 -16 7 -8
2 B1
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
44663 0
0
13 Logic Switch~
5 719 809 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21344 512
2 5V
-7 -16 7 -8
2 B2
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
44663 1
0
13 Logic Switch~
5 557 807 0 1 11
0 19
0
0 0 21344 512
2 0V
-7 -16 7 -8
2 B3
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
44663 2
0
13 Logic Switch~
5 409 806 0 1 11
0 21
0
0 0 21344 512
2 0V
-7 -16 7 -8
2 B4
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
44663 3
0
13 Logic Switch~
5 890 165 0 10 11
0 47 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
44663 4
0
13 Logic Switch~
5 713 168 0 1 11
0 48
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
44663 5
0
13 Logic Switch~
5 564 172 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
44663 6
0
13 Logic Switch~
5 429 172 0 1 11
0 50
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
44663 7
0
13 Logic Switch~
5 243 433 0 1 11
0 23
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4747 0 0
2
44663 8
0
13 Logic Switch~
5 175 435 0 1 11
0 22
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
44663 9
0
13 Logic Switch~
5 102 437 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
44663 10
0
13 Logic Switch~
5 95 532 0 1 11
0 11
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
44663 11
0
14 Logic Display~
6 1117 391 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
5 Carry
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
44663 12
0
14 Logic Display~
6 1142 389 0 1 2
10 36
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
44663 13
0
14 Logic Display~
6 1164 389 0 1 2
10 35
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
44663 14
0
14 Logic Display~
6 1188 387 0 1 2
10 34
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
44663 15
0
14 Logic Display~
6 1215 387 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
44663 16
0
9 Inverter~
13 111 480 0 2 22
0 13 12
0
0 0 608 270
6 74LS04
-21 -19 21 -11
3 NOT
20 -8 41 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 13 0
1 U
9323 0 0
2
44663 17
0
9 2-In AND~
219 365 523 0 3 22
0 12 11 10
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 12 0
1 U
317 0 0
2
44663 18
0
9 Inverter~
13 831 755 0 2 22
0 16 14
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 NOT
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 8 0
1 U
3108 0 0
2
44663 19
0
9 Inverter~
13 662 757 0 2 22
0 17 15
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 NOT
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 8 0
1 U
4299 0 0
2
44663 20
0
9 Inverter~
13 523 760 0 2 22
0 19 18
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 NOT
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 8 0
1 U
9672 0 0
2
44663 21
0
9 Inverter~
13 356 758 0 2 22
0 21 20
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 NOT
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 8 0
1 U
7876 0 0
2
44663 22
0
9 2-In AND~
219 860 613 0 3 22
0 23 16 25
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 11 0
1 U
6369 0 0
2
44663 23
0
9 2-In AND~
219 859 660 0 3 22
0 22 14 24
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 11 0
1 U
9172 0 0
2
44663 24
0
9 2-In AND~
219 692 620 0 3 22
0 23 17 27
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 11 0
1 U
7100 0 0
2
44663 25
0
9 2-In AND~
219 691 667 0 3 22
0 22 15 26
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
3820 0 0
2
44663 26
0
9 2-In AND~
219 551 623 0 3 22
0 23 19 29
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
7678 0 0
2
44663 27
0
9 2-In AND~
219 550 670 0 3 22
0 22 18 28
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
961 0 0
2
44663 28
0
9 2-In AND~
219 383 675 0 3 22
0 22 20 30
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
3178 0 0
2
44663 29
0
9 2-In AND~
219 384 628 0 3 22
0 23 21 31
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3409 0 0
2
44663 30
0
6 74LS83
105 1075 457 0 14 29
0 2 3 4 5 6 7 8 9 10
36 35 34 33 32
0
0 0 4832 0
5 74F83
-18 -60 17 -52
2 U1
-7 -61 7 -53
0
15 DVCC=5;DGND=12;
125 %D [%5bi %12bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%5bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 8 10 16 4 7 11 13
15 2 6 9 14 1 3 8 10 16
4 7 11 13 15 2 6 9 14 0
65 0 0 0 1 0 0 0
1 U
3951 0 0
2
44663 31
0
8 2-In OR~
219 907 572 0 3 22
0 25 24 9
0
0 0 608 90
6 74LS32
-21 -24 21 -16
2 OR
-3 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 9 0
1 U
8885 0 0
2
44663 32
0
8 2-In OR~
219 731 575 0 3 22
0 27 26 8
0
0 0 608 90
6 74LS32
-21 -24 21 -16
2 OR
-3 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 9 0
1 U
3780 0 0
2
44663 33
0
8 2-In OR~
219 582 578 0 3 22
0 29 28 7
0
0 0 608 90
6 74LS32
-21 -24 21 -16
2 OR
-3 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 9 0
1 U
9265 0 0
2
44663 34
0
8 2-In OR~
219 429 580 0 3 22
0 31 30 6
0
0 0 608 90
6 74LS32
-21 -24 21 -16
2 OR
-3 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 9 0
1 U
9442 0 0
2
44663 35
0
9 Inverter~
13 285 205 0 2 22
0 23 37
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 8 0
1 U
9424 0 0
2
44663 36
0
9 Inverter~
13 286 161 0 2 22
0 22 38
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 8 0
1 U
9968 0 0
2
44663 37
0
9 4-In AND~
219 869 208 0 5 22
0 13 38 37 16 44
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 AND
-15 -6 6 2
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 7 0
1 U
9281 0 0
2
44663 38
0
9 4-In AND~
219 868 258 0 5 22
0 13 22 37 14 43
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 AND
-13 -4 8 4
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 7 0
1 U
8464 0 0
2
44663 39
0
9 4-In AND~
219 696 216 0 5 22
0 13 38 37 17 46
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 AND
-15 -6 6 2
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 6 0
1 U
7168 0 0
2
44663 40
0
9 4-In AND~
219 695 267 0 5 22
0 13 22 37 15 45
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 6 0
1 U
3171 0 0
2
44663 41
0
9 4-In AND~
219 551 219 0 5 22
0 13 38 37 19 42
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 AND
-15 -6 6 2
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 5 0
1 U
4139 0 0
2
44663 42
0
9 4-In AND~
219 550 269 0 5 22
0 13 22 37 18 41
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 AND
-11 -4 10 4
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 5 0
1 U
6435 0 0
2
44663 43
0
9 4-In AND~
219 401 268 0 5 22
0 13 22 37 20 39
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 AND
-13 -5 8 3
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 12 13 8 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 2 4 0
1 U
5283 0 0
2
44663 44
0
9 4-In AND~
219 402 218 0 5 22
0 13 38 37 21 40
0
0 0 608 0
6 74LS21
-21 -28 21 -20
3 AND
-15 -6 6 2
0
15 DVCC=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 1 2 4 5 6 1 2 4 5
6 9 10 12 13 8 0 0 0 0
0 6 0
65 0 0 0 2 1 4 0
1 U
6874 0 0
2
44663 45
0
8 3-In OR~
219 907 350 0 4 22
0 47 44 43 5
0
0 0 608 270
4 4075
-14 -24 14 -16
2 OR
-2 1 12 9
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 3 0
1 U
5305 0 0
2
44663 46
0
8 3-In OR~
219 732 357 0 4 22
0 48 46 45 4
0
0 0 608 270
4 4075
-14 -24 14 -16
2 OR
-2 1 12 9
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 2 0
1 U
34 0 0
2
44663 47
0
8 3-In OR~
219 582 361 0 4 22
0 49 42 41 3
0
0 0 608 270
4 4075
-14 -24 14 -16
2 OR
-2 1 12 9
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 2 0
1 U
969 0 0
2
44663 48
0
8 3-In OR~
219 429 361 0 4 22
0 50 40 39 2
0
0 0 608 270
4 4075
-14 -24 14 -16
2 OR
-3 2 11 10
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 2 0
1 U
8402 0 0
2
44663 49
0
91
4 1 2 0 0 8320 0 50 32 0 0 3
432 391
432 421
1043 421
4 2 3 0 0 8320 0 49 32 0 0 3
585 391
585 430
1043 430
4 3 4 0 0 8320 0 48 32 0 0 3
735 387
735 439
1043 439
4 4 5 0 0 8320 0 47 32 0 0 3
910 380
910 448
1043 448
3 5 6 0 0 8320 0 36 32 0 0 3
432 550
432 457
1043 457
3 6 7 0 0 8320 0 35 32 0 0 3
585 548
585 466
1043 466
3 7 8 0 0 8320 0 34 32 0 0 3
734 545
734 475
1043 475
3 8 9 0 0 8320 0 33 32 0 0 3
910 542
910 484
1043 484
3 9 10 0 0 4224 0 19 32 0 0 4
386 523
1035 523
1035 502
1043 502
1 2 11 0 0 4224 0 12 19 0 0 2
107 532
341 532
2 1 12 0 0 8320 0 18 19 0 0 3
114 498
114 514
341 514
1 1 13 0 0 4096 0 11 18 0 0 2
114 437
114 462
0 4 14 0 0 8320 0 0 40 24 0 4
834 731
802 731
802 272
844 272
0 4 15 0 0 8320 0 0 42 25 0 4
665 732
631 732
631 281
671 281
4 0 16 0 0 8320 0 39 0 0 27 4
845 222
792 222
792 803
815 803
4 0 17 0 0 8320 0 41 0 0 28 4
672 230
622 230
622 809
651 809
4 0 18 0 0 8320 0 44 0 0 26 4
526 283
479 283
479 733
526 733
4 0 19 0 0 8320 0 43 0 0 29 4
527 233
471 233
471 807
511 807
4 0 20 0 0 8320 0 45 0 0 32 4
377 282
316 282
316 732
359 732
4 0 21 0 0 8320 0 46 0 0 31 4
378 232
308 232
308 806
344 806
1 0 19 0 0 0 0 22 0 0 29 2
526 778
526 807
1 0 17 0 0 0 0 21 0 0 28 2
665 775
665 809
1 0 16 0 0 0 0 20 0 0 27 2
834 773
834 803
2 2 14 0 0 0 0 25 20 0 0 3
835 669
834 669
834 737
2 2 15 0 0 0 0 27 21 0 0 3
667 676
665 676
665 739
2 2 18 0 0 0 0 29 22 0 0 2
526 679
526 742
2 1 16 0 0 0 0 24 1 0 0 4
836 622
815 622
815 803
886 803
2 1 17 0 0 0 0 26 2 0 0 4
668 629
651 629
651 809
707 809
2 1 19 0 0 0 0 28 3 0 0 4
527 632
511 632
511 807
545 807
1 0 21 0 0 0 0 23 0 0 31 2
359 776
359 806
1 2 21 0 0 0 0 4 31 0 0 4
397 806
344 806
344 637
360 637
2 2 20 0 0 0 0 23 30 0 0 2
359 740
359 684
1 0 22 0 0 8192 0 30 0 0 36 3
359 666
352 666
352 722
1 0 22 0 0 8192 0 29 0 0 36 3
526 661
517 661
517 722
1 0 22 0 0 8192 0 27 0 0 36 3
667 658
657 658
657 722
1 1 22 0 0 8320 0 10 25 0 0 5
187 435
187 722
824 722
824 651
835 651
1 0 23 0 0 8192 0 26 0 0 40 3
668 611
643 611
643 704
1 0 23 0 0 0 0 28 0 0 40 3
527 614
504 614
504 704
1 0 23 0 0 0 0 31 0 0 40 3
360 619
336 619
336 704
0 1 23 0 0 8320 0 0 24 59 0 6
262 433
262 704
807 704
807 605
836 605
836 604
3 2 24 0 0 8320 0 25 33 0 0 3
880 660
919 660
919 588
3 1 25 0 0 8320 0 24 33 0 0 3
881 613
901 613
901 588
3 2 26 0 0 8320 0 27 34 0 0 3
712 667
743 667
743 591
3 1 27 0 0 8320 0 26 34 0 0 3
713 620
725 620
725 591
3 2 28 0 0 8320 0 29 35 0 0 3
571 670
594 670
594 594
3 1 29 0 0 8320 0 28 35 0 0 3
572 623
576 623
576 594
3 2 30 0 0 8320 0 30 36 0 0 3
404 675
441 675
441 596
3 1 31 0 0 8320 0 31 36 0 0 3
405 628
423 628
423 596
14 1 32 0 0 8320 0 32 13 0 0 4
1107 502
1118 502
1118 409
1117 409
13 1 33 0 0 4224 0 32 17 0 0 3
1107 475
1215 475
1215 405
12 1 34 0 0 4224 0 32 16 0 0 3
1107 466
1188 466
1188 405
11 1 35 0 0 4224 0 32 15 0 0 3
1107 457
1164 457
1164 407
10 1 36 0 0 8320 0 32 14 0 0 3
1107 448
1142 448
1142 407
0 0 37 0 0 4096 0 0 0 57 74 2
320 205
320 273
0 0 22 0 0 0 0 0 0 60 75 2
187 176
329 176
0 0 13 0 0 4096 0 0 0 77 61 3
336 124
114 124
114 132
2 0 37 0 0 0 0 37 0 0 78 2
306 205
354 205
2 0 38 0 0 4096 0 38 0 0 79 2
307 161
364 161
1 1 23 0 0 0 0 9 37 0 0 4
255 433
262 433
262 205
270 205
1 1 22 0 0 0 0 10 38 0 0 3
187 435
187 161
271 161
1 0 13 0 0 4096 0 11 0 0 76 3
114 437
114 132
374 132
3 0 37 0 0 8192 0 42 0 0 74 3
671 272
630 272
630 57
2 0 22 0 0 0 0 42 0 0 75 3
671 263
638 263
638 66
1 0 13 0 0 0 0 42 0 0 77 3
671 254
645 254
645 74
3 0 37 0 0 8192 0 44 0 0 74 3
526 274
479 274
479 57
2 0 22 0 0 0 0 44 0 0 75 3
526 265
485 265
485 66
1 0 13 0 0 0 0 44 0 0 77 3
526 256
492 256
492 74
3 0 37 0 0 0 0 41 0 0 78 3
672 221
655 221
655 110
3 0 37 0 0 0 0 43 0 0 78 3
527 224
510 224
510 110
2 0 38 0 0 8192 0 41 0 0 79 3
672 212
661 212
661 121
2 0 38 0 0 8192 0 43 0 0 79 3
527 215
519 215
519 121
1 0 13 0 0 0 0 41 0 0 76 3
672 203
667 203
667 132
1 0 13 0 0 0 0 43 0 0 76 3
527 206
526 206
526 132
3 3 37 0 0 12416 0 45 40 0 0 6
377 273
320 273
320 57
804 57
804 263
844 263
2 2 22 0 0 0 0 45 40 0 0 6
377 264
329 264
329 66
812 66
812 254
844 254
1 1 13 0 0 12288 0 46 39 0 0 5
378 205
374 205
374 132
845 132
845 195
1 1 13 0 0 12416 0 45 40 0 0 6
377 255
336 255
336 74
819 74
819 245
844 245
3 3 37 0 0 0 0 46 39 0 0 6
378 223
354 223
354 110
829 110
829 213
845 213
2 2 38 0 0 12416 0 46 39 0 0 6
378 214
364 214
364 121
837 121
837 204
845 204
5 3 39 0 0 8320 0 45 50 0 0 3
422 268
423 268
423 345
5 2 40 0 0 8320 0 46 50 0 0 3
423 218
432 218
432 346
5 3 41 0 0 8320 0 44 49 0 0 3
571 269
576 269
576 345
5 2 42 0 0 8320 0 43 49 0 0 3
572 219
585 219
585 346
5 3 43 0 0 8320 0 40 47 0 0 3
889 258
901 258
901 334
5 2 44 0 0 8320 0 39 47 0 0 3
890 208
910 208
910 335
5 3 45 0 0 8320 0 42 48 0 0 3
716 267
726 267
726 341
5 2 46 0 0 8320 0 41 48 0 0 3
717 216
735 216
735 342
1 1 47 0 0 8320 0 5 47 0 0 3
902 165
919 165
919 334
1 1 48 0 0 8320 0 6 48 0 0 3
725 168
744 168
744 341
1 1 49 0 0 8320 0 7 49 0 0 3
576 172
594 172
594 345
1 1 50 0 0 4224 0 50 8 0 0 2
441 345
441 172
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
