CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 300 30 70 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
72
13 Logic Switch~
5 939 846 0 10 11
0 42 0 0 0 0 0 0 0 0
1
0
0 0 21344 512
2 5V
-7 -16 7 -8
2 B5
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.90027e-315 0
0
13 Logic Switch~
5 760 852 0 10 11
0 43 0 0 0 0 0 0 0 0
1
0
0 0 21344 512
2 5V
-7 -16 7 -8
2 B6
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.90027e-315 5.26354e-315
0
13 Logic Switch~
5 598 850 0 1 11
0 45
0
0 0 21344 512
2 0V
-7 -16 7 -8
2 B7
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.90027e-315 5.30499e-315
0
13 Logic Switch~
5 450 849 0 1 11
0 47
0
0 0 21344 512
2 0V
-7 -16 7 -8
2 B8
-7 -26 7 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.90027e-315 5.32571e-315
0
13 Logic Switch~
5 931 208 0 10 11
0 66 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.90027e-315 5.34643e-315
0
13 Logic Switch~
5 754 211 0 1 11
0 67
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5572 0 0
2
5.90027e-315 5.3568e-315
0
13 Logic Switch~
5 605 215 0 10 11
0 68 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 A3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.90027e-315 5.36716e-315
0
13 Logic Switch~
5 470 215 0 1 11
0 4
0
0 0 21344 0
2 0V
-6 -16 8 -8
2 A4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.90027e-315 5.37752e-315
0
13 Logic Switch~
5 284 476 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 S0
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.90027e-315 5.38788e-315
0
13 Logic Switch~
5 216 478 0 10 11
0 48 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 S1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
972 0 0
2
5.90027e-315 5.39306e-315
0
13 Logic Switch~
5 143 480 0 10 11
0 39 0 0 0 0 0 0 0 0
1
0
0 0 21344 0
2 5V
-6 -16 8 -8
2 S2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3472 0 0
2
5.90027e-315 5.39824e-315
0
13 Logic Switch~
5 136 575 0 1 11
0 38
0
0 0 21344 0
2 0V
-6 -16 8 -8
3 Cin
-9 -26 12 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9998 0 0
2
5.90027e-315 5.40342e-315
0
14 Logic Display~
6 1416 376 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
5 Carry
-17 -21 18 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.90027e-315 5.4086e-315
0
14 Logic Display~
6 1439 380 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4597 0 0
2
5.90027e-315 5.41378e-315
0
14 Logic Display~
6 1461 383 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
5.90027e-315 5.41896e-315
0
14 Logic Display~
6 1488 385 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.90027e-315 5.42414e-315
0
14 Logic Display~
6 1516 379 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
5.90027e-315 5.42933e-315
0
9 Inverter~
13 872 798 0 2 22
0 42 40
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 NOT
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 13 0
1 U
9323 0 0
2
5.90027e-315 5.43192e-315
0
9 Inverter~
13 703 800 0 2 22
0 43 41
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 NOT
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 13 0
1 U
317 0 0
2
5.90027e-315 5.43451e-315
0
9 Inverter~
13 564 803 0 2 22
0 45 44
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 NOT
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 13 0
1 U
3108 0 0
2
5.90027e-315 5.4371e-315
0
9 Inverter~
13 397 801 0 2 22
0 47 46
0
0 0 608 90
6 74LS04
-21 -19 21 -11
3 NOT
16 -2 37 6
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 13 0
1 U
4299 0 0
2
5.90027e-315 5.43969e-315
0
9 2-In AND~
219 901 656 0 3 22
0 49 42 51
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 12 0
1 U
9672 0 0
2
5.90027e-315 5.44228e-315
0
9 2-In AND~
219 900 703 0 3 22
0 48 40 50
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 12 0
1 U
7876 0 0
2
5.90027e-315 5.44487e-315
0
9 2-In AND~
219 733 663 0 3 22
0 49 43 53
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 14 0
1 U
6369 0 0
2
5.90027e-315 5.44746e-315
0
9 2-In AND~
219 732 710 0 3 22
0 48 41 52
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 14 0
1 U
9172 0 0
2
5.90027e-315 5.45005e-315
0
9 2-In AND~
219 592 666 0 3 22
0 49 45 55
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 14 0
1 U
7100 0 0
2
5.90027e-315 5.45264e-315
0
9 2-In AND~
219 591 713 0 3 22
0 48 44 54
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 14 0
1 U
3820 0 0
2
5.90027e-315 5.45523e-315
0
9 2-In AND~
219 424 718 0 3 22
0 48 46 56
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 15 0
1 U
7678 0 0
2
5.90027e-315 5.45782e-315
0
9 2-In AND~
219 425 671 0 3 22
0 49 47 57
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -6 7 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 15 0
1 U
961 0 0
2
5.90027e-315 5.46041e-315
0
8 2-In OR~
219 948 615 0 3 22
0 51 50 23
0
0 0 608 90
6 74LS32
-21 -24 21 -16
2 OR
-3 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 16 0
1 U
3178 0 0
2
5.90027e-315 5.463e-315
0
8 2-In OR~
219 772 618 0 3 22
0 53 52 36
0
0 0 608 90
6 74LS32
-21 -24 21 -16
2 OR
-3 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 16 0
1 U
3409 0 0
2
5.90027e-315 5.46559e-315
0
8 2-In OR~
219 623 621 0 3 22
0 55 54 31
0
0 0 608 90
6 74LS32
-21 -24 21 -16
2 OR
-3 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 16 0
1 U
3951 0 0
2
5.90027e-315 5.46818e-315
0
8 2-In OR~
219 470 623 0 3 22
0 57 56 27
0
0 0 608 90
6 74LS32
-21 -24 21 -16
2 OR
-3 -6 11 2
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 16 0
1 U
8885 0 0
2
5.90027e-315 5.47077e-315
0
9 Inverter~
13 326 248 0 2 22
0 49 58
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 17 0
1 U
3780 0 0
2
5.90027e-315 5.47207e-315
0
9 Inverter~
13 327 204 0 2 22
0 48 59
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 17 0
1 U
9265 0 0
2
5.90027e-315 5.47336e-315
0
8 3-In OR~
219 948 393 0 4 22
0 66 63 62 24
0
0 0 608 270
4 4075
-14 -24 14 -16
2 OR
-2 1 12 9
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 3 0
1 U
9442 0 0
2
5.90027e-315 5.47466e-315
0
8 3-In OR~
219 773 400 0 4 22
0 67 65 64 37
0
0 0 608 270
4 4075
-14 -24 14 -16
2 OR
-2 1 12 9
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 11 12 13 10 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 3 3 0
1 U
9424 0 0
2
5.90027e-315 5.47595e-315
0
8 3-In OR~
219 623 404 0 4 22
0 68 61 60 32
0
0 0 608 270
4 4075
-14 -24 14 -16
2 OR
-2 1 12 9
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 3 3 5 6 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 1 22 0
1 U
9968 0 0
2
5.90027e-315 5.47725e-315
0
8 3-In OR~
219 470 404 0 4 22
0 4 3 2 5
0
0 0 608 270
4 4075
-14 -24 14 -16
2 OR
-1 -1 13 7
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
17

0 1 2 8 9 3 3 5 6 1
2 8 9 11 12 13 10 0
65 0 0 0 3 2 22 0
1 U
9281 0 0
2
5.90027e-315 5.47854e-315
0
9 Inverter~
13 174 520 0 2 22
0 39 8
0
0 0 608 0
6 74LS04
-21 -19 21 -11
3 NOT
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 17 0
1 U
8464 0 0
2
5.90027e-315 5.47984e-315
0
9 2-In AND~
219 268 550 0 3 22
0 8 38 20
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 15 0
1 U
7168 0 0
2
5.90027e-315 5.48113e-315
0
5 4082~
219 444 261 0 5 22
0 39 59 58 47 3
0
0 0 608 0
4 4082
-7 -24 21 -16
3 AND
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 18 0
1 U
3171 0 0
2
5.90027e-315 5.48243e-315
0
5 4082~
219 441 311 0 5 22
0 39 48 58 46 2
0
0 0 608 0
4 4082
-7 -24 21 -16
3 AND
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 18 0
1 U
4139 0 0
2
5.90027e-315 5.48372e-315
0
5 4082~
219 739 259 0 5 22
0 39 59 58 43 65
0
0 0 608 0
4 4082
-7 -24 21 -16
3 AND
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 19 0
1 U
6435 0 0
2
5.90027e-315 5.48502e-315
0
5 4082~
219 594 262 0 5 22
0 39 59 58 45 61
0
0 0 608 0
4 4082
-7 -24 21 -16
3 AND
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 20 0
1 U
5283 0 0
2
5.90027e-315 5.48631e-315
0
5 4082~
219 591 312 0 5 22
0 39 48 58 44 60
0
0 0 608 0
4 4082
-7 -24 21 -16
3 AND
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 20 0
1 U
6874 0 0
2
5.90027e-315 5.48761e-315
0
5 4082~
219 737 310 0 5 22
0 39 48 58 41 64
0
0 0 608 0
4 4082
-7 -24 21 -16
3 AND
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 21 0
1 U
5305 0 0
2
5.90027e-315 5.4889e-315
0
5 4082~
219 910 251 0 5 22
0 39 59 58 42 63
0
0 0 608 0
4 4082
-7 -24 21 -16
3 AND
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 21 0
1 U
34 0 0
2
5.90027e-315 5.4902e-315
0
5 4082~
219 908 301 0 5 22
0 39 48 58 40 62
0
0 0 608 0
4 4082
-7 -24 21 -16
3 AND
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 23 0
1 U
969 0 0
2
5.90027e-315 5.49149e-315
0
8 2-In OR~
219 1282 716 0 3 22
0 35 34 11
0
0 0 608 0
6 74LS32
-21 -24 21 -16
2 OR
3 -5 17 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 31 0
1 U
8402 0 0
2
5.90027e-315 5.49279e-315
0
9 2-In AND~
219 1242 731 0 3 22
0 37 36 34
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -5 9 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 30 0
1 U
3751 0 0
2
5.90027e-315 5.49408e-315
0
9 2-In AND~
219 1242 694 0 3 22
0 13 9 35
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 30 0
1 U
4292 0 0
2
5.90027e-315 5.49538e-315
0
9 2-In XOR~
219 1277 659 0 3 22
0 13 9 18
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 XOR
-1 -5 20 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 29 0
1 U
6118 0 0
2
5.90027e-315 5.49667e-315
0
9 2-In XOR~
219 1177 638 0 3 22
0 37 36 13
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 XOR
-2 -5 19 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 29 0
1 U
34 0 0
2
5.90027e-315 5.49797e-315
0
9 2-In XOR~
219 1172 775 0 3 22
0 32 31 33
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 XOR
-2 -5 19 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 32 0
1 U
6357 0 0
2
5.90027e-315 5.49926e-315
0
9 2-In XOR~
219 1279 784 0 3 22
0 33 7 17
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 XOR
-1 -5 20 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 32 0
1 U
319 0 0
2
5.90027e-315 5.50056e-315
0
9 2-In AND~
219 1242 819 0 3 22
0 33 7 30
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 30 0
1 U
3976 0 0
2
5.90027e-315 5.50185e-315
0
9 2-In AND~
219 1241 857 0 3 22
0 32 31 29
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -5 9 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 33 0
1 U
7634 0 0
2
5.90027e-315 5.50315e-315
0
8 2-In OR~
219 1280 837 0 3 22
0 30 29 10
0
0 0 608 0
6 74LS32
-21 -24 21 -16
2 OR
3 -5 17 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 31 0
1 U
523 0 0
2
5.90027e-315 5.50444e-315
0
9 2-In XOR~
219 1174 902 0 3 22
0 5 27 28
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 XOR
-2 -5 19 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 9 10 8 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 32 0
1 U
6748 0 0
2
5.90027e-315 5.50574e-315
0
9 2-In XOR~
219 1279 911 0 3 22
0 28 6 16
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 XOR
-1 -5 20 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 32 0
1 U
6901 0 0
2
5.90027e-315 5.50703e-315
0
9 2-In AND~
219 1241 955 0 3 22
0 28 6 26
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 33 0
1 U
842 0 0
2
5.90027e-315 5.50833e-315
0
9 2-In AND~
219 1238 998 0 3 22
0 5 27 25
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -5 9 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 33 0
1 U
3277 0 0
2
5.90027e-315 5.50963e-315
0
8 2-In OR~
219 1282 980 0 3 22
0 26 25 15
0
0 0 608 0
6 74LS32
-21 -24 21 -16
2 OR
3 -5 17 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 31 0
1 U
4212 0 0
2
5.90027e-315 5.51092e-315
0
8 2-In OR~
219 1285 570 0 3 22
0 22 21 12
0
0 0 608 0
6 74LS32
-21 -24 21 -16
2 OR
3 -5 17 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 31 0
1 U
4720 0 0
2
5.90027e-315 5.51222e-315
0
9 2-In AND~
219 1241 589 0 3 22
0 24 23 21
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -5 9 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 30 0
1 U
5551 0 0
2
5.90027e-315 5.51286e-315
0
9 2-In AND~
219 1241 553 0 3 22
0 14 20 22
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-14 -4 7 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 28 0
1 U
6986 0 0
2
5.90027e-315 5.51351e-315
0
9 2-In XOR~
219 1277 509 0 3 22
0 14 20 19
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 XOR
-1 -5 20 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 29 0
1 U
8745 0 0
2
5.90027e-315 5.51416e-315
0
9 2-In XOR~
219 1178 489 0 3 22
0 24 23 14
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 XOR
0 -4 21 4
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 29 0
1 U
9592 0 0
2
5.90027e-315 5.51481e-315
0
9 2-In AND~
219 1339 579 0 3 22
0 12 8 9
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 33 0
1 U
8748 0 0
2
5.90027e-315 5.51545e-315
0
9 2-In AND~
219 1339 724 0 3 22
0 11 8 7
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 24 0
1 U
7168 0 0
2
5.90027e-315 5.5161e-315
0
9 2-In AND~
219 1336 845 0 3 22
0 10 8 6
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 25 0
1 U
631 0 0
2
5.90027e-315 5.51675e-315
0
128
5 3 2 0 0 8320 0 43 39 0 0 5
462 311
466 311
466 373
464 373
464 388
5 2 3 0 0 8320 0 42 39 0 0 3
465 261
473 261
473 389
1 1 4 0 0 4224 0 39 8 0 0 5
482 388
482 225
491 225
491 215
482 215
1 4 5 0 0 12416 0 60 39 0 0 5
1158 893
1003 893
1003 460
473 460
473 434
3 0 6 0 0 8320 0 72 0 0 14 5
1357 845
1357 880
1064 880
1064 940
1072 940
3 0 7 0 0 8320 0 71 0 0 15 5
1360 724
1360 760
1073 760
1073 813
1086 813
2 0 8 0 0 8192 0 72 0 0 9 3
1312 854
1312 870
980 870
2 0 8 0 0 8192 0 71 0 0 9 3
1315 733
1315 753
980 753
0 2 8 0 0 8320 0 0 70 55 0 6
201 520
201 870
980 870
980 609
1315 609
1315 588
0 3 9 0 0 12416 0 0 70 48 0 6
1084 689
1074 689
1074 619
1368 619
1368 579
1360 579
1 3 10 0 0 4224 0 72 59 0 0 3
1312 836
1312 837
1313 837
1 3 11 0 0 4224 0 71 50 0 0 2
1315 715
1315 716
1 3 12 0 0 4224 0 70 65 0 0 2
1315 570
1318 570
2 2 6 0 0 0 0 62 61 0 0 4
1217 964
1072 964
1072 920
1263 920
2 2 7 0 0 0 0 57 56 0 0 4
1218 828
1086 828
1086 793
1263 793
0 1 13 0 0 4224 0 0 52 17 0 3
1210 638
1210 685
1218 685
3 1 13 0 0 0 0 54 53 0 0 4
1210 638
1253 638
1253 650
1261 650
3 1 14 0 0 8320 0 69 67 0 0 4
1211 489
1212 489
1212 544
1217 544
3 1 15 0 0 8320 0 64 13 0 0 3
1315 980
1416 980
1416 394
3 1 16 0 0 8320 0 61 14 0 0 3
1312 911
1439 911
1439 398
3 1 17 0 0 8320 0 56 15 0 0 3
1312 784
1461 784
1461 401
3 1 18 0 0 8320 0 53 16 0 0 3
1310 659
1488 659
1488 403
3 1 19 0 0 4224 0 68 17 0 0 4
1310 509
1518 509
1518 397
1516 397
3 0 20 0 0 4224 0 41 0 0 29 2
289 550
1101 550
3 2 21 0 0 8320 0 66 65 0 0 4
1262 589
1267 589
1267 579
1272 579
3 1 22 0 0 8320 0 67 65 0 0 4
1262 553
1266 553
1266 561
1272 561
0 2 23 0 0 8192 0 0 66 30 0 3
1119 511
1119 598
1217 598
0 1 24 0 0 4096 0 0 66 32 0 3
1132 467
1132 580
1217 580
2 2 20 0 0 0 0 67 68 0 0 6
1217 562
1101 562
1101 531
1251 531
1251 518
1261 518
3 2 23 0 0 24704 0 30 69 0 0 9
951 585
951 528
1041 528
1041 526
1042 526
1042 511
1151 511
1151 498
1162 498
3 1 14 0 0 0 0 69 68 0 0 4
1211 489
1249 489
1249 500
1261 500
4 1 24 0 0 8320 0 36 69 0 0 7
951 423
951 491
1090 491
1090 467
1150 467
1150 480
1162 480
3 2 25 0 0 8320 0 63 64 0 0 4
1259 998
1263 998
1263 989
1269 989
3 1 26 0 0 8320 0 62 64 0 0 4
1262 955
1264 955
1264 971
1269 971
0 2 27 0 0 8192 0 0 63 38 0 3
1057 911
1057 1007
1214 1007
0 1 5 0 0 0 0 0 63 4 0 3
1087 893
1087 989
1214 989
1 0 28 0 0 8192 0 62 0 0 39 3
1217 946
1213 946
1213 902
3 2 27 0 0 8320 0 33 60 0 0 5
473 593
473 500
1011 500
1011 911
1158 911
3 1 28 0 0 4224 0 60 61 0 0 2
1207 902
1263 902
3 2 29 0 0 8320 0 58 59 0 0 4
1262 857
1265 857
1265 846
1267 846
3 1 30 0 0 8320 0 57 59 0 0 4
1263 819
1264 819
1264 828
1267 828
0 2 31 0 0 8192 0 0 58 45 0 3
1096 842
1096 866
1217 866
0 1 32 0 0 8192 0 0 58 47 0 3
1108 766
1108 848
1217 848
1 0 33 0 0 8192 0 57 0 0 46 3
1218 810
1205 810
1205 775
3 2 31 0 0 8320 0 32 55 0 0 7
626 591
626 509
1021 509
1021 842
1123 842
1123 784
1156 784
3 1 33 0 0 4224 0 55 56 0 0 2
1205 775
1263 775
4 1 32 0 0 8320 0 38 55 0 0 5
626 434
626 473
1066 473
1066 766
1156 766
2 2 9 0 0 0 0 52 53 0 0 4
1218 703
1084 703
1084 668
1261 668
3 2 34 0 0 8320 0 51 50 0 0 4
1263 731
1265 731
1265 725
1269 725
3 1 35 0 0 8320 0 52 50 0 0 4
1263 694
1265 694
1265 707
1269 707
0 2 36 0 0 8192 0 0 51 57 0 3
1096 647
1096 740
1218 740
0 1 37 0 0 8192 0 0 51 53 0 3
1109 629
1109 722
1218 722
4 1 37 0 0 8320 0 37 54 0 0 5
776 430
776 482
1080 482
1080 629
1161 629
1 2 38 0 0 4224 0 12 41 0 0 4
148 575
237 575
237 559
244 559
2 1 8 0 0 0 0 40 41 0 0 4
195 520
237 520
237 541
244 541
1 1 39 0 0 4096 0 11 40 0 0 3
155 480
155 520
159 520
3 2 36 0 0 8320 0 31 54 0 0 5
775 588
775 518
1033 518
1033 647
1161 647
0 4 40 0 0 8320 0 0 49 69 0 4
875 774
843 774
843 315
884 315
0 4 41 0 0 8320 0 0 47 70 0 4
706 775
672 775
672 324
713 324
4 0 42 0 0 8320 0 48 0 0 72 4
886 265
833 265
833 846
856 846
4 0 43 0 0 8320 0 44 0 0 73 4
715 273
663 273
663 852
692 852
4 0 44 0 0 8320 0 46 0 0 71 4
567 326
520 326
520 776
567 776
4 0 45 0 0 16512 0 45 0 0 74 6
570 276
572 276
572 276
512 276
512 850
552 850
4 0 46 0 0 8320 0 43 0 0 77 4
417 325
357 325
357 775
400 775
4 0 47 0 0 8320 0 42 0 0 76 4
420 275
349 275
349 849
385 849
1 0 45 0 0 0 0 20 0 0 74 2
567 821
567 850
1 0 43 0 0 0 0 19 0 0 73 2
706 818
706 852
1 0 42 0 0 0 0 18 0 0 72 2
875 816
875 846
2 2 40 0 0 0 0 23 18 0 0 3
876 712
875 712
875 780
2 2 41 0 0 0 0 25 19 0 0 3
708 719
706 719
706 782
2 2 44 0 0 0 0 27 20 0 0 2
567 722
567 785
2 1 42 0 0 0 0 22 1 0 0 4
877 665
856 665
856 846
927 846
2 1 43 0 0 0 0 24 2 0 0 4
709 672
692 672
692 852
748 852
2 1 45 0 0 0 0 26 3 0 0 4
568 675
552 675
552 850
586 850
1 0 47 0 0 0 0 21 0 0 76 2
400 819
400 849
1 2 47 0 0 0 0 4 29 0 0 4
438 849
385 849
385 680
401 680
2 2 46 0 0 0 0 21 28 0 0 2
400 783
400 727
1 0 48 0 0 8192 0 28 0 0 81 3
400 709
393 709
393 765
1 0 48 0 0 8192 0 27 0 0 81 3
567 704
558 704
558 765
1 0 48 0 0 8192 0 25 0 0 81 3
708 701
698 701
698 765
1 1 48 0 0 8320 0 10 23 0 0 5
228 478
228 765
865 765
865 694
876 694
1 0 49 0 0 8192 0 24 0 0 85 3
709 654
684 654
684 747
1 0 49 0 0 0 0 26 0 0 85 3
568 657
545 657
545 747
1 0 49 0 0 0 0 29 0 0 85 3
401 662
377 662
377 747
0 1 49 0 0 8320 0 0 22 99 0 5
303 476
303 747
848 747
848 647
877 647
3 2 50 0 0 8320 0 23 30 0 0 3
921 703
960 703
960 631
3 1 51 0 0 8320 0 22 30 0 0 3
922 656
942 656
942 631
3 2 52 0 0 8320 0 25 31 0 0 3
753 710
784 710
784 634
3 1 53 0 0 8320 0 24 31 0 0 3
754 663
766 663
766 634
3 2 54 0 0 8320 0 27 32 0 0 3
612 713
635 713
635 637
3 1 55 0 0 8320 0 26 32 0 0 3
613 666
617 666
617 637
3 2 56 0 0 8320 0 28 33 0 0 3
445 718
482 718
482 639
3 1 57 0 0 8320 0 29 33 0 0 3
446 671
464 671
464 639
0 0 58 0 0 4096 0 0 0 97 114 2
361 248
361 316
0 0 48 0 0 0 0 0 0 100 115 2
228 219
370 219
0 0 39 0 0 4096 0 0 0 117 101 3
377 167
155 167
155 175
2 0 58 0 0 0 0 34 0 0 118 2
347 248
395 248
2 0 59 0 0 4096 0 35 0 0 119 2
348 204
405 204
1 1 49 0 0 0 0 9 34 0 0 4
296 476
303 476
303 248
311 248
1 1 48 0 0 0 0 10 35 0 0 3
228 478
228 204
312 204
1 0 39 0 0 4096 0 11 0 0 116 3
155 480
155 175
415 175
3 0 58 0 0 8192 0 47 0 0 114 3
713 315
671 315
671 100
2 0 48 0 0 0 0 47 0 0 115 3
713 306
679 306
679 109
1 0 39 0 0 0 0 47 0 0 117 3
713 297
686 297
686 117
3 0 58 0 0 8192 0 46 0 0 114 3
567 317
520 317
520 100
2 0 48 0 0 0 0 46 0 0 115 3
567 308
526 308
526 109
1 0 39 0 0 0 0 46 0 0 117 3
567 299
533 299
533 117
3 0 58 0 0 0 0 44 0 0 118 3
715 264
696 264
696 153
3 0 58 0 0 0 0 45 0 0 118 5
570 267
572 267
572 267
551 267
551 153
2 0 59 0 0 8192 0 44 0 0 119 3
715 255
702 255
702 164
2 0 59 0 0 16384 0 45 0 0 119 5
570 258
572 258
572 258
560 258
560 164
1 0 39 0 0 0 0 44 0 0 116 3
715 246
708 246
708 175
1 0 39 0 0 0 0 45 0 0 116 5
570 249
572 249
572 249
567 249
567 175
3 3 58 0 0 12416 0 43 49 0 0 6
417 316
361 316
361 100
845 100
845 306
884 306
2 2 48 0 0 0 0 43 49 0 0 6
417 307
370 307
370 109
853 109
853 297
884 297
1 1 39 0 0 12288 0 42 48 0 0 5
420 248
415 248
415 175
886 175
886 238
1 1 39 0 0 12416 0 43 49 0 0 6
417 298
377 298
377 117
860 117
860 288
884 288
3 3 58 0 0 0 0 42 48 0 0 6
420 266
395 266
395 153
870 153
870 256
886 256
2 2 59 0 0 12416 0 42 48 0 0 6
420 257
405 257
405 164
878 164
878 247
886 247
5 3 60 0 0 8320 0 46 38 0 0 3
612 312
617 312
617 388
5 2 61 0 0 8320 0 45 38 0 0 3
615 262
626 262
626 389
5 3 62 0 0 8320 0 49 36 0 0 3
929 301
942 301
942 377
5 2 63 0 0 8320 0 48 36 0 0 3
931 251
951 251
951 378
5 3 64 0 0 8320 0 47 37 0 0 3
758 310
767 310
767 384
5 2 65 0 0 8320 0 44 37 0 0 3
760 259
776 259
776 385
1 1 66 0 0 8320 0 5 36 0 0 3
943 208
960 208
960 377
1 1 67 0 0 8320 0 6 37 0 0 3
766 211
785 211
785 384
1 1 68 0 0 8320 0 7 38 0 0 3
617 215
635 215
635 388
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
